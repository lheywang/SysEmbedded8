-- QsysTD.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity QsysTD is
	port (
		boutons_poussoirs_export : in  std_logic_vector(1 downto 0)  := (others => '0'); -- boutons_poussoirs.export
		clk_clk                  : in  std_logic                     := '0';             --               clk.clk
		hex1_export              : out std_logic_vector(31 downto 0);                    --              hex1.export
		hex2_export              : out std_logic_vector(31 downto 0);                    --              hex2.export
		interrupteurs_export     : in  std_logic_vector(9 downto 0)  := (others => '0'); --     interrupteurs.export
		leds_export              : out std_logic_vector(9 downto 0);                     --              leds.export
		pwm_ctrl_export          : out std_logic_vector(31 downto 0);                    --          pwm_ctrl.export
		pwm_status_export        : in  std_logic_vector(7 downto 0)  := (others => '0'); --        pwm_status.export
		reset_reset_n            : in  std_logic                     := '0'              --             reset.reset_n
	);
end entity QsysTD;

architecture rtl of QsysTD is
	component QsysTD_BOUTONS_POUSSOIRS is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component QsysTD_BOUTONS_POUSSOIRS;

	component QsysTD_HEX3_HEX0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component QsysTD_HEX3_HEX0;

	component QsysTD_INTERRUPTEURS is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(9 downto 0)  := (others => 'X')  -- export
		);
	end component QsysTD_INTERRUPTEURS;

	component QsysTD_LEDR is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(9 downto 0)                      -- export
		);
	end component QsysTD_LEDR;

	component QsysTD_MEMOIRE_ONCHIP is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component QsysTD_MEMOIRE_ONCHIP;

	component QsysTD_NiosII_CPU is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(18 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(18 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component QsysTD_NiosII_CPU;

	component QsysTD_PWM_CTRL is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(31 downto 0)                     -- export
		);
	end component QsysTD_PWM_CTRL;

	component QsysTD_PWM_STATUS is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component QsysTD_PWM_STATUS;

	component QsysTD_SYS_CLK_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component QsysTD_SYS_CLK_timer;

	component QsysTD_SYS_MEL is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component QsysTD_SYS_MEL;

	component QsysTD_SYS_SEC is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component QsysTD_SYS_SEC;

	component QsysTD_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component QsysTD_jtag_uart_0;

	component QsysTD_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component QsysTD_sysid_qsys_0;

	component QsysTD_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                 : in  std_logic                     := 'X';             -- clk
			jtag_uart_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			NiosII_CPU_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			NiosII_CPU_data_master_address                : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			NiosII_CPU_data_master_waitrequest            : out std_logic;                                        -- waitrequest
			NiosII_CPU_data_master_byteenable             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			NiosII_CPU_data_master_read                   : in  std_logic                     := 'X';             -- read
			NiosII_CPU_data_master_readdata               : out std_logic_vector(31 downto 0);                    -- readdata
			NiosII_CPU_data_master_write                  : in  std_logic                     := 'X';             -- write
			NiosII_CPU_data_master_writedata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			NiosII_CPU_data_master_debugaccess            : in  std_logic                     := 'X';             -- debugaccess
			NiosII_CPU_instruction_master_address         : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			NiosII_CPU_instruction_master_waitrequest     : out std_logic;                                        -- waitrequest
			NiosII_CPU_instruction_master_read            : in  std_logic                     := 'X';             -- read
			NiosII_CPU_instruction_master_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			NiosII_CPU_instruction_master_readdatavalid   : out std_logic;                                        -- readdatavalid
			BOUTONS_POUSSOIRS_s1_address                  : out std_logic_vector(1 downto 0);                     -- address
			BOUTONS_POUSSOIRS_s1_write                    : out std_logic;                                        -- write
			BOUTONS_POUSSOIRS_s1_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			BOUTONS_POUSSOIRS_s1_writedata                : out std_logic_vector(31 downto 0);                    -- writedata
			BOUTONS_POUSSOIRS_s1_chipselect               : out std_logic;                                        -- chipselect
			HEX3_HEX0_s1_address                          : out std_logic_vector(1 downto 0);                     -- address
			HEX3_HEX0_s1_write                            : out std_logic;                                        -- write
			HEX3_HEX0_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			HEX3_HEX0_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			HEX3_HEX0_s1_chipselect                       : out std_logic;                                        -- chipselect
			HEX5_HEX4_s1_address                          : out std_logic_vector(1 downto 0);                     -- address
			HEX5_HEX4_s1_write                            : out std_logic;                                        -- write
			HEX5_HEX4_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			HEX5_HEX4_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			HEX5_HEX4_s1_chipselect                       : out std_logic;                                        -- chipselect
			INTERRUPTEURS_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			INTERRUPTEURS_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_address         : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write           : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read            : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata       : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest     : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect      : out std_logic;                                        -- chipselect
			LEDR_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			LEDR_s1_write                                 : out std_logic;                                        -- write
			LEDR_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			LEDR_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			LEDR_s1_chipselect                            : out std_logic;                                        -- chipselect
			MEMOIRE_ONCHIP_s1_address                     : out std_logic_vector(14 downto 0);                    -- address
			MEMOIRE_ONCHIP_s1_write                       : out std_logic;                                        -- write
			MEMOIRE_ONCHIP_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			MEMOIRE_ONCHIP_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			MEMOIRE_ONCHIP_s1_byteenable                  : out std_logic_vector(3 downto 0);                     -- byteenable
			MEMOIRE_ONCHIP_s1_chipselect                  : out std_logic;                                        -- chipselect
			MEMOIRE_ONCHIP_s1_clken                       : out std_logic;                                        -- clken
			NiosII_CPU_debug_mem_slave_address            : out std_logic_vector(8 downto 0);                     -- address
			NiosII_CPU_debug_mem_slave_write              : out std_logic;                                        -- write
			NiosII_CPU_debug_mem_slave_read               : out std_logic;                                        -- read
			NiosII_CPU_debug_mem_slave_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			NiosII_CPU_debug_mem_slave_writedata          : out std_logic_vector(31 downto 0);                    -- writedata
			NiosII_CPU_debug_mem_slave_byteenable         : out std_logic_vector(3 downto 0);                     -- byteenable
			NiosII_CPU_debug_mem_slave_waitrequest        : in  std_logic                     := 'X';             -- waitrequest
			NiosII_CPU_debug_mem_slave_debugaccess        : out std_logic;                                        -- debugaccess
			PWM_CTRL_s1_address                           : out std_logic_vector(1 downto 0);                     -- address
			PWM_CTRL_s1_write                             : out std_logic;                                        -- write
			PWM_CTRL_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PWM_CTRL_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			PWM_CTRL_s1_chipselect                        : out std_logic;                                        -- chipselect
			PWM_STATUS_s1_address                         : out std_logic_vector(1 downto 0);                     -- address
			PWM_STATUS_s1_write                           : out std_logic;                                        -- write
			PWM_STATUS_s1_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PWM_STATUS_s1_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			PWM_STATUS_s1_chipselect                      : out std_logic;                                        -- chipselect
			SYS_CLK_timer_s1_address                      : out std_logic_vector(2 downto 0);                     -- address
			SYS_CLK_timer_s1_write                        : out std_logic;                                        -- write
			SYS_CLK_timer_s1_readdata                     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SYS_CLK_timer_s1_writedata                    : out std_logic_vector(15 downto 0);                    -- writedata
			SYS_CLK_timer_s1_chipselect                   : out std_logic;                                        -- chipselect
			SYS_MEL_s1_address                            : out std_logic_vector(2 downto 0);                     -- address
			SYS_MEL_s1_write                              : out std_logic;                                        -- write
			SYS_MEL_s1_readdata                           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SYS_MEL_s1_writedata                          : out std_logic_vector(15 downto 0);                    -- writedata
			SYS_MEL_s1_chipselect                         : out std_logic;                                        -- chipselect
			SYS_SEC_s1_address                            : out std_logic_vector(2 downto 0);                     -- address
			SYS_SEC_s1_write                              : out std_logic;                                        -- write
			SYS_SEC_s1_readdata                           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SYS_SEC_s1_writedata                          : out std_logic_vector(15 downto 0);                    -- writedata
			SYS_SEC_s1_chipselect                         : out std_logic;                                        -- chipselect
			sysid_qsys_0_control_slave_address            : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata           : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component QsysTD_mm_interconnect_0;

	component QsysTD_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			receiver5_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component QsysTD_irq_mapper;

	component qsystd_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component qsystd_rst_controller;

	component qsystd_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component qsystd_rst_controller_001;

	signal niosii_cpu_data_master_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:NiosII_CPU_data_master_readdata -> NiosII_CPU:d_readdata
	signal niosii_cpu_data_master_waitrequest                              : std_logic;                     -- mm_interconnect_0:NiosII_CPU_data_master_waitrequest -> NiosII_CPU:d_waitrequest
	signal niosii_cpu_data_master_debugaccess                              : std_logic;                     -- NiosII_CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NiosII_CPU_data_master_debugaccess
	signal niosii_cpu_data_master_address                                  : std_logic_vector(18 downto 0); -- NiosII_CPU:d_address -> mm_interconnect_0:NiosII_CPU_data_master_address
	signal niosii_cpu_data_master_byteenable                               : std_logic_vector(3 downto 0);  -- NiosII_CPU:d_byteenable -> mm_interconnect_0:NiosII_CPU_data_master_byteenable
	signal niosii_cpu_data_master_read                                     : std_logic;                     -- NiosII_CPU:d_read -> mm_interconnect_0:NiosII_CPU_data_master_read
	signal niosii_cpu_data_master_write                                    : std_logic;                     -- NiosII_CPU:d_write -> mm_interconnect_0:NiosII_CPU_data_master_write
	signal niosii_cpu_data_master_writedata                                : std_logic_vector(31 downto 0); -- NiosII_CPU:d_writedata -> mm_interconnect_0:NiosII_CPU_data_master_writedata
	signal niosii_cpu_instruction_master_readdata                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:NiosII_CPU_instruction_master_readdata -> NiosII_CPU:i_readdata
	signal niosii_cpu_instruction_master_waitrequest                       : std_logic;                     -- mm_interconnect_0:NiosII_CPU_instruction_master_waitrequest -> NiosII_CPU:i_waitrequest
	signal niosii_cpu_instruction_master_address                           : std_logic_vector(18 downto 0); -- NiosII_CPU:i_address -> mm_interconnect_0:NiosII_CPU_instruction_master_address
	signal niosii_cpu_instruction_master_read                              : std_logic;                     -- NiosII_CPU:i_read -> mm_interconnect_0:NiosII_CPU_instruction_master_read
	signal niosii_cpu_instruction_master_readdatavalid                     : std_logic;                     -- mm_interconnect_0:NiosII_CPU_instruction_master_readdatavalid -> NiosII_CPU:i_readdatavalid
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata           : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address            : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_niosii_cpu_debug_mem_slave_readdata           : std_logic_vector(31 downto 0); -- NiosII_CPU:debug_mem_slave_readdata -> mm_interconnect_0:NiosII_CPU_debug_mem_slave_readdata
	signal mm_interconnect_0_niosii_cpu_debug_mem_slave_waitrequest        : std_logic;                     -- NiosII_CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:NiosII_CPU_debug_mem_slave_waitrequest
	signal mm_interconnect_0_niosii_cpu_debug_mem_slave_debugaccess        : std_logic;                     -- mm_interconnect_0:NiosII_CPU_debug_mem_slave_debugaccess -> NiosII_CPU:debug_mem_slave_debugaccess
	signal mm_interconnect_0_niosii_cpu_debug_mem_slave_address            : std_logic_vector(8 downto 0);  -- mm_interconnect_0:NiosII_CPU_debug_mem_slave_address -> NiosII_CPU:debug_mem_slave_address
	signal mm_interconnect_0_niosii_cpu_debug_mem_slave_read               : std_logic;                     -- mm_interconnect_0:NiosII_CPU_debug_mem_slave_read -> NiosII_CPU:debug_mem_slave_read
	signal mm_interconnect_0_niosii_cpu_debug_mem_slave_byteenable         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:NiosII_CPU_debug_mem_slave_byteenable -> NiosII_CPU:debug_mem_slave_byteenable
	signal mm_interconnect_0_niosii_cpu_debug_mem_slave_write              : std_logic;                     -- mm_interconnect_0:NiosII_CPU_debug_mem_slave_write -> NiosII_CPU:debug_mem_slave_write
	signal mm_interconnect_0_niosii_cpu_debug_mem_slave_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:NiosII_CPU_debug_mem_slave_writedata -> NiosII_CPU:debug_mem_slave_writedata
	signal mm_interconnect_0_memoire_onchip_s1_chipselect                  : std_logic;                     -- mm_interconnect_0:MEMOIRE_ONCHIP_s1_chipselect -> MEMOIRE_ONCHIP:chipselect
	signal mm_interconnect_0_memoire_onchip_s1_readdata                    : std_logic_vector(31 downto 0); -- MEMOIRE_ONCHIP:readdata -> mm_interconnect_0:MEMOIRE_ONCHIP_s1_readdata
	signal mm_interconnect_0_memoire_onchip_s1_address                     : std_logic_vector(14 downto 0); -- mm_interconnect_0:MEMOIRE_ONCHIP_s1_address -> MEMOIRE_ONCHIP:address
	signal mm_interconnect_0_memoire_onchip_s1_byteenable                  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:MEMOIRE_ONCHIP_s1_byteenable -> MEMOIRE_ONCHIP:byteenable
	signal mm_interconnect_0_memoire_onchip_s1_write                       : std_logic;                     -- mm_interconnect_0:MEMOIRE_ONCHIP_s1_write -> MEMOIRE_ONCHIP:write
	signal mm_interconnect_0_memoire_onchip_s1_writedata                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:MEMOIRE_ONCHIP_s1_writedata -> MEMOIRE_ONCHIP:writedata
	signal mm_interconnect_0_memoire_onchip_s1_clken                       : std_logic;                     -- mm_interconnect_0:MEMOIRE_ONCHIP_s1_clken -> MEMOIRE_ONCHIP:clken
	signal mm_interconnect_0_sys_clk_timer_s1_chipselect                   : std_logic;                     -- mm_interconnect_0:SYS_CLK_timer_s1_chipselect -> SYS_CLK_timer:chipselect
	signal mm_interconnect_0_sys_clk_timer_s1_readdata                     : std_logic_vector(15 downto 0); -- SYS_CLK_timer:readdata -> mm_interconnect_0:SYS_CLK_timer_s1_readdata
	signal mm_interconnect_0_sys_clk_timer_s1_address                      : std_logic_vector(2 downto 0);  -- mm_interconnect_0:SYS_CLK_timer_s1_address -> SYS_CLK_timer:address
	signal mm_interconnect_0_sys_clk_timer_s1_write                        : std_logic;                     -- mm_interconnect_0:SYS_CLK_timer_s1_write -> mm_interconnect_0_sys_clk_timer_s1_write:in
	signal mm_interconnect_0_sys_clk_timer_s1_writedata                    : std_logic_vector(15 downto 0); -- mm_interconnect_0:SYS_CLK_timer_s1_writedata -> SYS_CLK_timer:writedata
	signal mm_interconnect_0_interrupteurs_s1_readdata                     : std_logic_vector(31 downto 0); -- INTERRUPTEURS:readdata -> mm_interconnect_0:INTERRUPTEURS_s1_readdata
	signal mm_interconnect_0_interrupteurs_s1_address                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:INTERRUPTEURS_s1_address -> INTERRUPTEURS:address
	signal mm_interconnect_0_hex3_hex0_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:HEX3_HEX0_s1_chipselect -> HEX3_HEX0:chipselect
	signal mm_interconnect_0_hex3_hex0_s1_readdata                         : std_logic_vector(31 downto 0); -- HEX3_HEX0:readdata -> mm_interconnect_0:HEX3_HEX0_s1_readdata
	signal mm_interconnect_0_hex3_hex0_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:HEX3_HEX0_s1_address -> HEX3_HEX0:address
	signal mm_interconnect_0_hex3_hex0_s1_write                            : std_logic;                     -- mm_interconnect_0:HEX3_HEX0_s1_write -> mm_interconnect_0_hex3_hex0_s1_write:in
	signal mm_interconnect_0_hex3_hex0_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:HEX3_HEX0_s1_writedata -> HEX3_HEX0:writedata
	signal mm_interconnect_0_hex5_hex4_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:HEX5_HEX4_s1_chipselect -> HEX5_HEX4:chipselect
	signal mm_interconnect_0_hex5_hex4_s1_readdata                         : std_logic_vector(31 downto 0); -- HEX5_HEX4:readdata -> mm_interconnect_0:HEX5_HEX4_s1_readdata
	signal mm_interconnect_0_hex5_hex4_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:HEX5_HEX4_s1_address -> HEX5_HEX4:address
	signal mm_interconnect_0_hex5_hex4_s1_write                            : std_logic;                     -- mm_interconnect_0:HEX5_HEX4_s1_write -> mm_interconnect_0_hex5_hex4_s1_write:in
	signal mm_interconnect_0_hex5_hex4_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:HEX5_HEX4_s1_writedata -> HEX5_HEX4:writedata
	signal mm_interconnect_0_pwm_ctrl_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:PWM_CTRL_s1_chipselect -> PWM_CTRL:chipselect
	signal mm_interconnect_0_pwm_ctrl_s1_readdata                          : std_logic_vector(31 downto 0); -- PWM_CTRL:readdata -> mm_interconnect_0:PWM_CTRL_s1_readdata
	signal mm_interconnect_0_pwm_ctrl_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:PWM_CTRL_s1_address -> PWM_CTRL:address
	signal mm_interconnect_0_pwm_ctrl_s1_write                             : std_logic;                     -- mm_interconnect_0:PWM_CTRL_s1_write -> mm_interconnect_0_pwm_ctrl_s1_write:in
	signal mm_interconnect_0_pwm_ctrl_s1_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:PWM_CTRL_s1_writedata -> PWM_CTRL:writedata
	signal mm_interconnect_0_sys_sec_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:SYS_SEC_s1_chipselect -> SYS_SEC:chipselect
	signal mm_interconnect_0_sys_sec_s1_readdata                           : std_logic_vector(15 downto 0); -- SYS_SEC:readdata -> mm_interconnect_0:SYS_SEC_s1_readdata
	signal mm_interconnect_0_sys_sec_s1_address                            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:SYS_SEC_s1_address -> SYS_SEC:address
	signal mm_interconnect_0_sys_sec_s1_write                              : std_logic;                     -- mm_interconnect_0:SYS_SEC_s1_write -> mm_interconnect_0_sys_sec_s1_write:in
	signal mm_interconnect_0_sys_sec_s1_writedata                          : std_logic_vector(15 downto 0); -- mm_interconnect_0:SYS_SEC_s1_writedata -> SYS_SEC:writedata
	signal mm_interconnect_0_sys_mel_s1_chipselect                         : std_logic;                     -- mm_interconnect_0:SYS_MEL_s1_chipselect -> SYS_MEL:chipselect
	signal mm_interconnect_0_sys_mel_s1_readdata                           : std_logic_vector(15 downto 0); -- SYS_MEL:readdata -> mm_interconnect_0:SYS_MEL_s1_readdata
	signal mm_interconnect_0_sys_mel_s1_address                            : std_logic_vector(2 downto 0);  -- mm_interconnect_0:SYS_MEL_s1_address -> SYS_MEL:address
	signal mm_interconnect_0_sys_mel_s1_write                              : std_logic;                     -- mm_interconnect_0:SYS_MEL_s1_write -> mm_interconnect_0_sys_mel_s1_write:in
	signal mm_interconnect_0_sys_mel_s1_writedata                          : std_logic_vector(15 downto 0); -- mm_interconnect_0:SYS_MEL_s1_writedata -> SYS_MEL:writedata
	signal mm_interconnect_0_boutons_poussoirs_s1_chipselect               : std_logic;                     -- mm_interconnect_0:BOUTONS_POUSSOIRS_s1_chipselect -> BOUTONS_POUSSOIRS:chipselect
	signal mm_interconnect_0_boutons_poussoirs_s1_readdata                 : std_logic_vector(31 downto 0); -- BOUTONS_POUSSOIRS:readdata -> mm_interconnect_0:BOUTONS_POUSSOIRS_s1_readdata
	signal mm_interconnect_0_boutons_poussoirs_s1_address                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:BOUTONS_POUSSOIRS_s1_address -> BOUTONS_POUSSOIRS:address
	signal mm_interconnect_0_boutons_poussoirs_s1_write                    : std_logic;                     -- mm_interconnect_0:BOUTONS_POUSSOIRS_s1_write -> mm_interconnect_0_boutons_poussoirs_s1_write:in
	signal mm_interconnect_0_boutons_poussoirs_s1_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:BOUTONS_POUSSOIRS_s1_writedata -> BOUTONS_POUSSOIRS:writedata
	signal mm_interconnect_0_pwm_status_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:PWM_STATUS_s1_chipselect -> PWM_STATUS:chipselect
	signal mm_interconnect_0_pwm_status_s1_readdata                        : std_logic_vector(31 downto 0); -- PWM_STATUS:readdata -> mm_interconnect_0:PWM_STATUS_s1_readdata
	signal mm_interconnect_0_pwm_status_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:PWM_STATUS_s1_address -> PWM_STATUS:address
	signal mm_interconnect_0_pwm_status_s1_write                           : std_logic;                     -- mm_interconnect_0:PWM_STATUS_s1_write -> mm_interconnect_0_pwm_status_s1_write:in
	signal mm_interconnect_0_pwm_status_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:PWM_STATUS_s1_writedata -> PWM_STATUS:writedata
	signal mm_interconnect_0_ledr_s1_chipselect                            : std_logic;                     -- mm_interconnect_0:LEDR_s1_chipselect -> LEDR:chipselect
	signal mm_interconnect_0_ledr_s1_readdata                              : std_logic_vector(31 downto 0); -- LEDR:readdata -> mm_interconnect_0:LEDR_s1_readdata
	signal mm_interconnect_0_ledr_s1_address                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:LEDR_s1_address -> LEDR:address
	signal mm_interconnect_0_ledr_s1_write                                 : std_logic;                     -- mm_interconnect_0:LEDR_s1_write -> mm_interconnect_0_ledr_s1_write:in
	signal mm_interconnect_0_ledr_s1_writedata                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:LEDR_s1_writedata -> LEDR:writedata
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                        : std_logic;                     -- SYS_CLK_timer:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                        : std_logic;                     -- SYS_SEC:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                        : std_logic;                     -- SYS_MEL:irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                        : std_logic;                     -- BOUTONS_POUSSOIRS:irq -> irq_mapper:receiver4_irq
	signal irq_mapper_receiver5_irq                                        : std_logic;                     -- PWM_STATUS:irq -> irq_mapper:receiver5_irq
	signal niosii_cpu_irq_irq                                              : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> NiosII_CPU:irq
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset                              : std_logic;                     -- rst_controller_001:reset_out -> [MEMOIRE_ONCHIP:reset, irq_mapper:reset, mm_interconnect_0:NiosII_CPU_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset_req                          : std_logic;                     -- rst_controller_001:reset_req -> [MEMOIRE_ONCHIP:reset_req, NiosII_CPU:reset_req, rst_translator:reset_req_in]
	signal niosii_cpu_debug_reset_request_reset                            : std_logic;                     -- NiosII_CPU:debug_reset_request -> rst_controller_001:reset_in1
	signal reset_reset_n_ports_inv                                         : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_sys_clk_timer_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_0_sys_clk_timer_s1_write:inv -> SYS_CLK_timer:write_n
	signal mm_interconnect_0_hex3_hex0_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_hex3_hex0_s1_write:inv -> HEX3_HEX0:write_n
	signal mm_interconnect_0_hex5_hex4_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_hex5_hex4_s1_write:inv -> HEX5_HEX4:write_n
	signal mm_interconnect_0_pwm_ctrl_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_pwm_ctrl_s1_write:inv -> PWM_CTRL:write_n
	signal mm_interconnect_0_sys_sec_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_sys_sec_s1_write:inv -> SYS_SEC:write_n
	signal mm_interconnect_0_sys_mel_s1_write_ports_inv                    : std_logic;                     -- mm_interconnect_0_sys_mel_s1_write:inv -> SYS_MEL:write_n
	signal mm_interconnect_0_boutons_poussoirs_s1_write_ports_inv          : std_logic;                     -- mm_interconnect_0_boutons_poussoirs_s1_write:inv -> BOUTONS_POUSSOIRS:write_n
	signal mm_interconnect_0_pwm_status_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_pwm_status_s1_write:inv -> PWM_STATUS:write_n
	signal mm_interconnect_0_ledr_s1_write_ports_inv                       : std_logic;                     -- mm_interconnect_0_ledr_s1_write:inv -> LEDR:write_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> [BOUTONS_POUSSOIRS:reset_n, HEX3_HEX0:reset_n, HEX5_HEX4:reset_n, INTERRUPTEURS:reset_n, LEDR:reset_n, PWM_CTRL:reset_n, PWM_STATUS:reset_n, SYS_CLK_timer:reset_n, SYS_MEL:reset_n, SYS_SEC:reset_n, jtag_uart_0:rst_n, sysid_qsys_0:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                    : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> NiosII_CPU:reset_n

begin

	boutons_poussoirs : component QsysTD_BOUTONS_POUSSOIRS
		port map (
			clk        => clk_clk,                                                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,               --               reset.reset_n
			address    => mm_interconnect_0_boutons_poussoirs_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_boutons_poussoirs_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_boutons_poussoirs_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_boutons_poussoirs_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_boutons_poussoirs_s1_readdata,        --                    .readdata
			in_port    => boutons_poussoirs_export,                               -- external_connection.export
			irq        => irq_mapper_receiver4_irq                                --                 irq.irq
		);

	hex3_hex0 : component QsysTD_HEX3_HEX0
		port map (
			clk        => clk_clk,                                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_hex3_hex0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex3_hex0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex3_hex0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex3_hex0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex3_hex0_s1_readdata,        --                    .readdata
			out_port   => hex1_export                                     -- external_connection.export
		);

	hex5_hex4 : component QsysTD_HEX3_HEX0
		port map (
			clk        => clk_clk,                                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_hex5_hex4_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex5_hex4_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex5_hex4_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex5_hex4_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex5_hex4_s1_readdata,        --                    .readdata
			out_port   => hex2_export                                     -- external_connection.export
		);

	interrupteurs : component QsysTD_INTERRUPTEURS
		port map (
			clk      => clk_clk,                                     --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address  => mm_interconnect_0_interrupteurs_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_interrupteurs_s1_readdata, --                    .readdata
			in_port  => interrupteurs_export                         -- external_connection.export
		);

	ledr : component QsysTD_LEDR
		port map (
			clk        => clk_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_ledr_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_ledr_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_ledr_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_ledr_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_ledr_s1_readdata,        --                    .readdata
			out_port   => leds_export                                -- external_connection.export
		);

	memoire_onchip : component QsysTD_MEMOIRE_ONCHIP
		port map (
			clk        => clk_clk,                                        --   clk1.clk
			address    => mm_interconnect_0_memoire_onchip_s1_address,    --     s1.address
			clken      => mm_interconnect_0_memoire_onchip_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_memoire_onchip_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_memoire_onchip_s1_write,      --       .write
			readdata   => mm_interconnect_0_memoire_onchip_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_memoire_onchip_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_memoire_onchip_s1_byteenable, --       .byteenable
			reset      => rst_controller_001_reset_out_reset,             -- reset1.reset
			reset_req  => rst_controller_001_reset_out_reset_req,         --       .reset_req
			freeze     => '0'                                             -- (terminated)
		);

	niosii_cpu : component QsysTD_NiosII_CPU
		port map (
			clk                                 => clk_clk,                                                  --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,             --                     reset.reset_n
			reset_req                           => rst_controller_001_reset_out_reset_req,                   --                          .reset_req
			d_address                           => niosii_cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => niosii_cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => niosii_cpu_data_master_read,                              --                          .read
			d_readdata                          => niosii_cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => niosii_cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => niosii_cpu_data_master_write,                             --                          .write
			d_writedata                         => niosii_cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => niosii_cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => niosii_cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => niosii_cpu_instruction_master_read,                       --                          .read
			i_readdata                          => niosii_cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => niosii_cpu_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => niosii_cpu_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => niosii_cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => niosii_cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_niosii_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_niosii_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_niosii_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_niosii_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_niosii_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_niosii_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_niosii_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_niosii_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                      -- custom_instruction_master.readra
		);

	pwm_ctrl : component QsysTD_PWM_CTRL
		port map (
			clk        => clk_clk,                                       --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_pwm_ctrl_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pwm_ctrl_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pwm_ctrl_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pwm_ctrl_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pwm_ctrl_s1_readdata,        --                    .readdata
			out_port   => pwm_ctrl_export                                -- external_connection.export
		);

	pwm_status : component QsysTD_PWM_STATUS
		port map (
			clk        => clk_clk,                                         --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_0_pwm_status_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pwm_status_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pwm_status_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pwm_status_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pwm_status_s1_readdata,        --                    .readdata
			in_port    => pwm_status_export,                               -- external_connection.export
			irq        => irq_mapper_receiver5_irq                         --                 irq.irq
		);

	sys_clk_timer : component QsysTD_SYS_CLK_timer
		port map (
			clk        => clk_clk,                                            --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           -- reset.reset_n
			address    => mm_interconnect_0_sys_clk_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_sys_clk_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_sys_clk_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_sys_clk_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_sys_clk_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                            --   irq.irq
		);

	sys_mel : component QsysTD_SYS_MEL
		port map (
			clk        => clk_clk,                                      --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_sys_mel_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_sys_mel_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_sys_mel_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_sys_mel_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_sys_mel_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver3_irq                      --   irq.irq
		);

	sys_sec : component QsysTD_SYS_SEC
		port map (
			clk        => clk_clk,                                      --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_sys_sec_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_sys_sec_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_sys_sec_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_sys_sec_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_sys_sec_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver2_irq                      --   irq.irq
		);

	jtag_uart_0 : component QsysTD_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                         --               irq.irq
		);

	sysid_qsys_0 : component QsysTD_sysid_qsys_0
		port map (
			clock    => clk_clk,                                                 --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component QsysTD_mm_interconnect_0
		port map (
			clk_0_clk_clk                                 => clk_clk,                                                     --                               clk_0_clk.clk
			jtag_uart_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                              -- jtag_uart_0_reset_reset_bridge_in_reset.reset
			NiosII_CPU_reset_reset_bridge_in_reset_reset  => rst_controller_001_reset_out_reset,                          --  NiosII_CPU_reset_reset_bridge_in_reset.reset
			NiosII_CPU_data_master_address                => niosii_cpu_data_master_address,                              --                  NiosII_CPU_data_master.address
			NiosII_CPU_data_master_waitrequest            => niosii_cpu_data_master_waitrequest,                          --                                        .waitrequest
			NiosII_CPU_data_master_byteenable             => niosii_cpu_data_master_byteenable,                           --                                        .byteenable
			NiosII_CPU_data_master_read                   => niosii_cpu_data_master_read,                                 --                                        .read
			NiosII_CPU_data_master_readdata               => niosii_cpu_data_master_readdata,                             --                                        .readdata
			NiosII_CPU_data_master_write                  => niosii_cpu_data_master_write,                                --                                        .write
			NiosII_CPU_data_master_writedata              => niosii_cpu_data_master_writedata,                            --                                        .writedata
			NiosII_CPU_data_master_debugaccess            => niosii_cpu_data_master_debugaccess,                          --                                        .debugaccess
			NiosII_CPU_instruction_master_address         => niosii_cpu_instruction_master_address,                       --           NiosII_CPU_instruction_master.address
			NiosII_CPU_instruction_master_waitrequest     => niosii_cpu_instruction_master_waitrequest,                   --                                        .waitrequest
			NiosII_CPU_instruction_master_read            => niosii_cpu_instruction_master_read,                          --                                        .read
			NiosII_CPU_instruction_master_readdata        => niosii_cpu_instruction_master_readdata,                      --                                        .readdata
			NiosII_CPU_instruction_master_readdatavalid   => niosii_cpu_instruction_master_readdatavalid,                 --                                        .readdatavalid
			BOUTONS_POUSSOIRS_s1_address                  => mm_interconnect_0_boutons_poussoirs_s1_address,              --                    BOUTONS_POUSSOIRS_s1.address
			BOUTONS_POUSSOIRS_s1_write                    => mm_interconnect_0_boutons_poussoirs_s1_write,                --                                        .write
			BOUTONS_POUSSOIRS_s1_readdata                 => mm_interconnect_0_boutons_poussoirs_s1_readdata,             --                                        .readdata
			BOUTONS_POUSSOIRS_s1_writedata                => mm_interconnect_0_boutons_poussoirs_s1_writedata,            --                                        .writedata
			BOUTONS_POUSSOIRS_s1_chipselect               => mm_interconnect_0_boutons_poussoirs_s1_chipselect,           --                                        .chipselect
			HEX3_HEX0_s1_address                          => mm_interconnect_0_hex3_hex0_s1_address,                      --                            HEX3_HEX0_s1.address
			HEX3_HEX0_s1_write                            => mm_interconnect_0_hex3_hex0_s1_write,                        --                                        .write
			HEX3_HEX0_s1_readdata                         => mm_interconnect_0_hex3_hex0_s1_readdata,                     --                                        .readdata
			HEX3_HEX0_s1_writedata                        => mm_interconnect_0_hex3_hex0_s1_writedata,                    --                                        .writedata
			HEX3_HEX0_s1_chipselect                       => mm_interconnect_0_hex3_hex0_s1_chipselect,                   --                                        .chipselect
			HEX5_HEX4_s1_address                          => mm_interconnect_0_hex5_hex4_s1_address,                      --                            HEX5_HEX4_s1.address
			HEX5_HEX4_s1_write                            => mm_interconnect_0_hex5_hex4_s1_write,                        --                                        .write
			HEX5_HEX4_s1_readdata                         => mm_interconnect_0_hex5_hex4_s1_readdata,                     --                                        .readdata
			HEX5_HEX4_s1_writedata                        => mm_interconnect_0_hex5_hex4_s1_writedata,                    --                                        .writedata
			HEX5_HEX4_s1_chipselect                       => mm_interconnect_0_hex5_hex4_s1_chipselect,                   --                                        .chipselect
			INTERRUPTEURS_s1_address                      => mm_interconnect_0_interrupteurs_s1_address,                  --                        INTERRUPTEURS_s1.address
			INTERRUPTEURS_s1_readdata                     => mm_interconnect_0_interrupteurs_s1_readdata,                 --                                        .readdata
			jtag_uart_0_avalon_jtag_slave_address         => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,     --           jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write           => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,       --                                        .write
			jtag_uart_0_avalon_jtag_slave_read            => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,        --                                        .read
			jtag_uart_0_avalon_jtag_slave_readdata        => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,    --                                        .readdata
			jtag_uart_0_avalon_jtag_slave_writedata       => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,   --                                        .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest, --                                        .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,  --                                        .chipselect
			LEDR_s1_address                               => mm_interconnect_0_ledr_s1_address,                           --                                 LEDR_s1.address
			LEDR_s1_write                                 => mm_interconnect_0_ledr_s1_write,                             --                                        .write
			LEDR_s1_readdata                              => mm_interconnect_0_ledr_s1_readdata,                          --                                        .readdata
			LEDR_s1_writedata                             => mm_interconnect_0_ledr_s1_writedata,                         --                                        .writedata
			LEDR_s1_chipselect                            => mm_interconnect_0_ledr_s1_chipselect,                        --                                        .chipselect
			MEMOIRE_ONCHIP_s1_address                     => mm_interconnect_0_memoire_onchip_s1_address,                 --                       MEMOIRE_ONCHIP_s1.address
			MEMOIRE_ONCHIP_s1_write                       => mm_interconnect_0_memoire_onchip_s1_write,                   --                                        .write
			MEMOIRE_ONCHIP_s1_readdata                    => mm_interconnect_0_memoire_onchip_s1_readdata,                --                                        .readdata
			MEMOIRE_ONCHIP_s1_writedata                   => mm_interconnect_0_memoire_onchip_s1_writedata,               --                                        .writedata
			MEMOIRE_ONCHIP_s1_byteenable                  => mm_interconnect_0_memoire_onchip_s1_byteenable,              --                                        .byteenable
			MEMOIRE_ONCHIP_s1_chipselect                  => mm_interconnect_0_memoire_onchip_s1_chipselect,              --                                        .chipselect
			MEMOIRE_ONCHIP_s1_clken                       => mm_interconnect_0_memoire_onchip_s1_clken,                   --                                        .clken
			NiosII_CPU_debug_mem_slave_address            => mm_interconnect_0_niosii_cpu_debug_mem_slave_address,        --              NiosII_CPU_debug_mem_slave.address
			NiosII_CPU_debug_mem_slave_write              => mm_interconnect_0_niosii_cpu_debug_mem_slave_write,          --                                        .write
			NiosII_CPU_debug_mem_slave_read               => mm_interconnect_0_niosii_cpu_debug_mem_slave_read,           --                                        .read
			NiosII_CPU_debug_mem_slave_readdata           => mm_interconnect_0_niosii_cpu_debug_mem_slave_readdata,       --                                        .readdata
			NiosII_CPU_debug_mem_slave_writedata          => mm_interconnect_0_niosii_cpu_debug_mem_slave_writedata,      --                                        .writedata
			NiosII_CPU_debug_mem_slave_byteenable         => mm_interconnect_0_niosii_cpu_debug_mem_slave_byteenable,     --                                        .byteenable
			NiosII_CPU_debug_mem_slave_waitrequest        => mm_interconnect_0_niosii_cpu_debug_mem_slave_waitrequest,    --                                        .waitrequest
			NiosII_CPU_debug_mem_slave_debugaccess        => mm_interconnect_0_niosii_cpu_debug_mem_slave_debugaccess,    --                                        .debugaccess
			PWM_CTRL_s1_address                           => mm_interconnect_0_pwm_ctrl_s1_address,                       --                             PWM_CTRL_s1.address
			PWM_CTRL_s1_write                             => mm_interconnect_0_pwm_ctrl_s1_write,                         --                                        .write
			PWM_CTRL_s1_readdata                          => mm_interconnect_0_pwm_ctrl_s1_readdata,                      --                                        .readdata
			PWM_CTRL_s1_writedata                         => mm_interconnect_0_pwm_ctrl_s1_writedata,                     --                                        .writedata
			PWM_CTRL_s1_chipselect                        => mm_interconnect_0_pwm_ctrl_s1_chipselect,                    --                                        .chipselect
			PWM_STATUS_s1_address                         => mm_interconnect_0_pwm_status_s1_address,                     --                           PWM_STATUS_s1.address
			PWM_STATUS_s1_write                           => mm_interconnect_0_pwm_status_s1_write,                       --                                        .write
			PWM_STATUS_s1_readdata                        => mm_interconnect_0_pwm_status_s1_readdata,                    --                                        .readdata
			PWM_STATUS_s1_writedata                       => mm_interconnect_0_pwm_status_s1_writedata,                   --                                        .writedata
			PWM_STATUS_s1_chipselect                      => mm_interconnect_0_pwm_status_s1_chipselect,                  --                                        .chipselect
			SYS_CLK_timer_s1_address                      => mm_interconnect_0_sys_clk_timer_s1_address,                  --                        SYS_CLK_timer_s1.address
			SYS_CLK_timer_s1_write                        => mm_interconnect_0_sys_clk_timer_s1_write,                    --                                        .write
			SYS_CLK_timer_s1_readdata                     => mm_interconnect_0_sys_clk_timer_s1_readdata,                 --                                        .readdata
			SYS_CLK_timer_s1_writedata                    => mm_interconnect_0_sys_clk_timer_s1_writedata,                --                                        .writedata
			SYS_CLK_timer_s1_chipselect                   => mm_interconnect_0_sys_clk_timer_s1_chipselect,               --                                        .chipselect
			SYS_MEL_s1_address                            => mm_interconnect_0_sys_mel_s1_address,                        --                              SYS_MEL_s1.address
			SYS_MEL_s1_write                              => mm_interconnect_0_sys_mel_s1_write,                          --                                        .write
			SYS_MEL_s1_readdata                           => mm_interconnect_0_sys_mel_s1_readdata,                       --                                        .readdata
			SYS_MEL_s1_writedata                          => mm_interconnect_0_sys_mel_s1_writedata,                      --                                        .writedata
			SYS_MEL_s1_chipselect                         => mm_interconnect_0_sys_mel_s1_chipselect,                     --                                        .chipselect
			SYS_SEC_s1_address                            => mm_interconnect_0_sys_sec_s1_address,                        --                              SYS_SEC_s1.address
			SYS_SEC_s1_write                              => mm_interconnect_0_sys_sec_s1_write,                          --                                        .write
			SYS_SEC_s1_readdata                           => mm_interconnect_0_sys_sec_s1_readdata,                       --                                        .readdata
			SYS_SEC_s1_writedata                          => mm_interconnect_0_sys_sec_s1_writedata,                      --                                        .writedata
			SYS_SEC_s1_chipselect                         => mm_interconnect_0_sys_sec_s1_chipselect,                     --                                        .chipselect
			sysid_qsys_0_control_slave_address            => mm_interconnect_0_sysid_qsys_0_control_slave_address,        --              sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata           => mm_interconnect_0_sysid_qsys_0_control_slave_readdata        --                                        .readdata
		);

	irq_mapper : component QsysTD_irq_mapper
		port map (
			clk           => clk_clk,                            --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,           -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,           -- receiver4.irq
			receiver5_irq => irq_mapper_receiver5_irq,           -- receiver5.irq
			sender_irq    => niosii_cpu_irq_irq                  --    sender.irq
		);

	rst_controller : component qsystd_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component qsystd_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => niosii_cpu_debug_reset_request_reset,   -- reset_in1.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_sys_clk_timer_s1_write_ports_inv <= not mm_interconnect_0_sys_clk_timer_s1_write;

	mm_interconnect_0_hex3_hex0_s1_write_ports_inv <= not mm_interconnect_0_hex3_hex0_s1_write;

	mm_interconnect_0_hex5_hex4_s1_write_ports_inv <= not mm_interconnect_0_hex5_hex4_s1_write;

	mm_interconnect_0_pwm_ctrl_s1_write_ports_inv <= not mm_interconnect_0_pwm_ctrl_s1_write;

	mm_interconnect_0_sys_sec_s1_write_ports_inv <= not mm_interconnect_0_sys_sec_s1_write;

	mm_interconnect_0_sys_mel_s1_write_ports_inv <= not mm_interconnect_0_sys_mel_s1_write;

	mm_interconnect_0_boutons_poussoirs_s1_write_ports_inv <= not mm_interconnect_0_boutons_poussoirs_s1_write;

	mm_interconnect_0_pwm_status_s1_write_ports_inv <= not mm_interconnect_0_pwm_status_s1_write;

	mm_interconnect_0_ledr_s1_write_ports_inv <= not mm_interconnect_0_ledr_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of QsysTD
