// QsysTD.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module QsysTD (
		input  wire [1:0]  boutons_poussoirs_export, // boutons_poussoirs.export
		input  wire        clk_clk,                  //               clk.clk
		output wire [31:0] hex1_export,              //              hex1.export
		output wire [31:0] hex2_export,              //              hex2.export
		input  wire [9:0]  interrupteurs_export,     //     interrupteurs.export
		output wire [9:0]  leds_export,              //              leds.export
		output wire [31:0] pwm_ctrl_export,          //          pwm_ctrl.export
		input  wire [7:0]  pwm_status_export,        //        pwm_status.export
		input  wire        reset_reset_n             //             reset.reset_n
	);

	wire  [31:0] niosii_cpu_data_master_readdata;                             // mm_interconnect_0:NiosII_CPU_data_master_readdata -> NiosII_CPU:d_readdata
	wire         niosii_cpu_data_master_waitrequest;                          // mm_interconnect_0:NiosII_CPU_data_master_waitrequest -> NiosII_CPU:d_waitrequest
	wire         niosii_cpu_data_master_debugaccess;                          // NiosII_CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NiosII_CPU_data_master_debugaccess
	wire  [18:0] niosii_cpu_data_master_address;                              // NiosII_CPU:d_address -> mm_interconnect_0:NiosII_CPU_data_master_address
	wire   [3:0] niosii_cpu_data_master_byteenable;                           // NiosII_CPU:d_byteenable -> mm_interconnect_0:NiosII_CPU_data_master_byteenable
	wire         niosii_cpu_data_master_read;                                 // NiosII_CPU:d_read -> mm_interconnect_0:NiosII_CPU_data_master_read
	wire         niosii_cpu_data_master_write;                                // NiosII_CPU:d_write -> mm_interconnect_0:NiosII_CPU_data_master_write
	wire  [31:0] niosii_cpu_data_master_writedata;                            // NiosII_CPU:d_writedata -> mm_interconnect_0:NiosII_CPU_data_master_writedata
	wire  [31:0] niosii_cpu_instruction_master_readdata;                      // mm_interconnect_0:NiosII_CPU_instruction_master_readdata -> NiosII_CPU:i_readdata
	wire         niosii_cpu_instruction_master_waitrequest;                   // mm_interconnect_0:NiosII_CPU_instruction_master_waitrequest -> NiosII_CPU:i_waitrequest
	wire  [18:0] niosii_cpu_instruction_master_address;                       // NiosII_CPU:i_address -> mm_interconnect_0:NiosII_CPU_instruction_master_address
	wire         niosii_cpu_instruction_master_read;                          // NiosII_CPU:i_read -> mm_interconnect_0:NiosII_CPU_instruction_master_read
	wire         niosii_cpu_instruction_master_readdatavalid;                 // mm_interconnect_0:NiosII_CPU_instruction_master_readdatavalid -> NiosII_CPU:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_niosii_cpu_debug_mem_slave_readdata;       // NiosII_CPU:debug_mem_slave_readdata -> mm_interconnect_0:NiosII_CPU_debug_mem_slave_readdata
	wire         mm_interconnect_0_niosii_cpu_debug_mem_slave_waitrequest;    // NiosII_CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:NiosII_CPU_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_niosii_cpu_debug_mem_slave_debugaccess;    // mm_interconnect_0:NiosII_CPU_debug_mem_slave_debugaccess -> NiosII_CPU:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_niosii_cpu_debug_mem_slave_address;        // mm_interconnect_0:NiosII_CPU_debug_mem_slave_address -> NiosII_CPU:debug_mem_slave_address
	wire         mm_interconnect_0_niosii_cpu_debug_mem_slave_read;           // mm_interconnect_0:NiosII_CPU_debug_mem_slave_read -> NiosII_CPU:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_niosii_cpu_debug_mem_slave_byteenable;     // mm_interconnect_0:NiosII_CPU_debug_mem_slave_byteenable -> NiosII_CPU:debug_mem_slave_byteenable
	wire         mm_interconnect_0_niosii_cpu_debug_mem_slave_write;          // mm_interconnect_0:NiosII_CPU_debug_mem_slave_write -> NiosII_CPU:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_niosii_cpu_debug_mem_slave_writedata;      // mm_interconnect_0:NiosII_CPU_debug_mem_slave_writedata -> NiosII_CPU:debug_mem_slave_writedata
	wire         mm_interconnect_0_memoire_onchip_s1_chipselect;              // mm_interconnect_0:MEMOIRE_ONCHIP_s1_chipselect -> MEMOIRE_ONCHIP:chipselect
	wire  [31:0] mm_interconnect_0_memoire_onchip_s1_readdata;                // MEMOIRE_ONCHIP:readdata -> mm_interconnect_0:MEMOIRE_ONCHIP_s1_readdata
	wire  [14:0] mm_interconnect_0_memoire_onchip_s1_address;                 // mm_interconnect_0:MEMOIRE_ONCHIP_s1_address -> MEMOIRE_ONCHIP:address
	wire   [3:0] mm_interconnect_0_memoire_onchip_s1_byteenable;              // mm_interconnect_0:MEMOIRE_ONCHIP_s1_byteenable -> MEMOIRE_ONCHIP:byteenable
	wire         mm_interconnect_0_memoire_onchip_s1_write;                   // mm_interconnect_0:MEMOIRE_ONCHIP_s1_write -> MEMOIRE_ONCHIP:write
	wire  [31:0] mm_interconnect_0_memoire_onchip_s1_writedata;               // mm_interconnect_0:MEMOIRE_ONCHIP_s1_writedata -> MEMOIRE_ONCHIP:writedata
	wire         mm_interconnect_0_memoire_onchip_s1_clken;                   // mm_interconnect_0:MEMOIRE_ONCHIP_s1_clken -> MEMOIRE_ONCHIP:clken
	wire         mm_interconnect_0_sys_clk_timer_s1_chipselect;               // mm_interconnect_0:SYS_CLK_timer_s1_chipselect -> SYS_CLK_timer:chipselect
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_readdata;                 // SYS_CLK_timer:readdata -> mm_interconnect_0:SYS_CLK_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_clk_timer_s1_address;                  // mm_interconnect_0:SYS_CLK_timer_s1_address -> SYS_CLK_timer:address
	wire         mm_interconnect_0_sys_clk_timer_s1_write;                    // mm_interconnect_0:SYS_CLK_timer_s1_write -> SYS_CLK_timer:write_n
	wire  [15:0] mm_interconnect_0_sys_clk_timer_s1_writedata;                // mm_interconnect_0:SYS_CLK_timer_s1_writedata -> SYS_CLK_timer:writedata
	wire  [31:0] mm_interconnect_0_interrupteurs_s1_readdata;                 // INTERRUPTEURS:readdata -> mm_interconnect_0:INTERRUPTEURS_s1_readdata
	wire   [1:0] mm_interconnect_0_interrupteurs_s1_address;                  // mm_interconnect_0:INTERRUPTEURS_s1_address -> INTERRUPTEURS:address
	wire         mm_interconnect_0_ledr_s1_chipselect;                        // mm_interconnect_0:LEDR_s1_chipselect -> LEDR:chipselect
	wire  [31:0] mm_interconnect_0_ledr_s1_readdata;                          // LEDR:readdata -> mm_interconnect_0:LEDR_s1_readdata
	wire   [1:0] mm_interconnect_0_ledr_s1_address;                           // mm_interconnect_0:LEDR_s1_address -> LEDR:address
	wire         mm_interconnect_0_ledr_s1_write;                             // mm_interconnect_0:LEDR_s1_write -> LEDR:write_n
	wire  [31:0] mm_interconnect_0_ledr_s1_writedata;                         // mm_interconnect_0:LEDR_s1_writedata -> LEDR:writedata
	wire         mm_interconnect_0_hex3_hex0_s1_chipselect;                   // mm_interconnect_0:HEX3_HEX0_s1_chipselect -> HEX3_HEX0:chipselect
	wire  [31:0] mm_interconnect_0_hex3_hex0_s1_readdata;                     // HEX3_HEX0:readdata -> mm_interconnect_0:HEX3_HEX0_s1_readdata
	wire   [1:0] mm_interconnect_0_hex3_hex0_s1_address;                      // mm_interconnect_0:HEX3_HEX0_s1_address -> HEX3_HEX0:address
	wire         mm_interconnect_0_hex3_hex0_s1_write;                        // mm_interconnect_0:HEX3_HEX0_s1_write -> HEX3_HEX0:write_n
	wire  [31:0] mm_interconnect_0_hex3_hex0_s1_writedata;                    // mm_interconnect_0:HEX3_HEX0_s1_writedata -> HEX3_HEX0:writedata
	wire         mm_interconnect_0_hex5_hex4_s1_chipselect;                   // mm_interconnect_0:HEX5_HEX4_s1_chipselect -> HEX5_HEX4:chipselect
	wire  [31:0] mm_interconnect_0_hex5_hex4_s1_readdata;                     // HEX5_HEX4:readdata -> mm_interconnect_0:HEX5_HEX4_s1_readdata
	wire   [1:0] mm_interconnect_0_hex5_hex4_s1_address;                      // mm_interconnect_0:HEX5_HEX4_s1_address -> HEX5_HEX4:address
	wire         mm_interconnect_0_hex5_hex4_s1_write;                        // mm_interconnect_0:HEX5_HEX4_s1_write -> HEX5_HEX4:write_n
	wire  [31:0] mm_interconnect_0_hex5_hex4_s1_writedata;                    // mm_interconnect_0:HEX5_HEX4_s1_writedata -> HEX5_HEX4:writedata
	wire         mm_interconnect_0_pwm_ctrl_s1_chipselect;                    // mm_interconnect_0:PWM_CTRL_s1_chipselect -> PWM_CTRL:chipselect
	wire  [31:0] mm_interconnect_0_pwm_ctrl_s1_readdata;                      // PWM_CTRL:readdata -> mm_interconnect_0:PWM_CTRL_s1_readdata
	wire   [1:0] mm_interconnect_0_pwm_ctrl_s1_address;                       // mm_interconnect_0:PWM_CTRL_s1_address -> PWM_CTRL:address
	wire         mm_interconnect_0_pwm_ctrl_s1_write;                         // mm_interconnect_0:PWM_CTRL_s1_write -> PWM_CTRL:write_n
	wire  [31:0] mm_interconnect_0_pwm_ctrl_s1_writedata;                     // mm_interconnect_0:PWM_CTRL_s1_writedata -> PWM_CTRL:writedata
	wire         mm_interconnect_0_sys_sec_s1_chipselect;                     // mm_interconnect_0:SYS_SEC_s1_chipselect -> SYS_SEC:chipselect
	wire  [15:0] mm_interconnect_0_sys_sec_s1_readdata;                       // SYS_SEC:readdata -> mm_interconnect_0:SYS_SEC_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_sec_s1_address;                        // mm_interconnect_0:SYS_SEC_s1_address -> SYS_SEC:address
	wire         mm_interconnect_0_sys_sec_s1_write;                          // mm_interconnect_0:SYS_SEC_s1_write -> SYS_SEC:write_n
	wire  [15:0] mm_interconnect_0_sys_sec_s1_writedata;                      // mm_interconnect_0:SYS_SEC_s1_writedata -> SYS_SEC:writedata
	wire         mm_interconnect_0_sys_mel_s1_chipselect;                     // mm_interconnect_0:SYS_MEL_s1_chipselect -> SYS_MEL:chipselect
	wire  [15:0] mm_interconnect_0_sys_mel_s1_readdata;                       // SYS_MEL:readdata -> mm_interconnect_0:SYS_MEL_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_mel_s1_address;                        // mm_interconnect_0:SYS_MEL_s1_address -> SYS_MEL:address
	wire         mm_interconnect_0_sys_mel_s1_write;                          // mm_interconnect_0:SYS_MEL_s1_write -> SYS_MEL:write_n
	wire  [15:0] mm_interconnect_0_sys_mel_s1_writedata;                      // mm_interconnect_0:SYS_MEL_s1_writedata -> SYS_MEL:writedata
	wire         mm_interconnect_0_boutons_poussoirs_s1_chipselect;           // mm_interconnect_0:BOUTONS_POUSSOIRS_s1_chipselect -> BOUTONS_POUSSOIRS:chipselect
	wire  [31:0] mm_interconnect_0_boutons_poussoirs_s1_readdata;             // BOUTONS_POUSSOIRS:readdata -> mm_interconnect_0:BOUTONS_POUSSOIRS_s1_readdata
	wire   [1:0] mm_interconnect_0_boutons_poussoirs_s1_address;              // mm_interconnect_0:BOUTONS_POUSSOIRS_s1_address -> BOUTONS_POUSSOIRS:address
	wire         mm_interconnect_0_boutons_poussoirs_s1_write;                // mm_interconnect_0:BOUTONS_POUSSOIRS_s1_write -> BOUTONS_POUSSOIRS:write_n
	wire  [31:0] mm_interconnect_0_boutons_poussoirs_s1_writedata;            // mm_interconnect_0:BOUTONS_POUSSOIRS_s1_writedata -> BOUTONS_POUSSOIRS:writedata
	wire         mm_interconnect_0_pwm_status_s1_chipselect;                  // mm_interconnect_0:PWM_STATUS_s1_chipselect -> PWM_STATUS:chipselect
	wire  [31:0] mm_interconnect_0_pwm_status_s1_readdata;                    // PWM_STATUS:readdata -> mm_interconnect_0:PWM_STATUS_s1_readdata
	wire   [1:0] mm_interconnect_0_pwm_status_s1_address;                     // mm_interconnect_0:PWM_STATUS_s1_address -> PWM_STATUS:address
	wire         mm_interconnect_0_pwm_status_s1_write;                       // mm_interconnect_0:PWM_STATUS_s1_write -> PWM_STATUS:write_n
	wire  [31:0] mm_interconnect_0_pwm_status_s1_writedata;                   // mm_interconnect_0:PWM_STATUS_s1_writedata -> PWM_STATUS:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // SYS_CLK_timer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // SYS_SEC:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                    // SYS_MEL:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                    // BOUTONS_POUSSOIRS:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                    // PWM_STATUS:irq -> irq_mapper:receiver5_irq
	wire  [31:0] niosii_cpu_irq_irq;                                          // irq_mapper:sender_irq -> NiosII_CPU:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [BOUTONS_POUSSOIRS:reset_n, HEX3_HEX0:reset_n, HEX5_HEX4:reset_n, INTERRUPTEURS:reset_n, LEDR:reset_n, PWM_CTRL:reset_n, PWM_STATUS:reset_n, SYS_CLK_timer:reset_n, SYS_MEL:reset_n, SYS_SEC:reset_n, jtag_uart_0:rst_n, mm_interconnect_0:jtag_uart_0_reset_reset_bridge_in_reset_reset, sysid_qsys_0:reset_n]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [MEMOIRE_ONCHIP:reset, NiosII_CPU:reset_n, irq_mapper:reset, mm_interconnect_0:NiosII_CPU_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [MEMOIRE_ONCHIP:reset_req, NiosII_CPU:reset_req, rst_translator:reset_req_in]
	wire         niosii_cpu_debug_reset_request_reset;                        // NiosII_CPU:debug_reset_request -> rst_controller_001:reset_in1

	QsysTD_BOUTONS_POUSSOIRS boutons_poussoirs (
		.clk        (clk_clk),                                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_boutons_poussoirs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_boutons_poussoirs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_boutons_poussoirs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_boutons_poussoirs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_boutons_poussoirs_s1_readdata),   //                    .readdata
		.in_port    (boutons_poussoirs_export),                          // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                           //                 irq.irq
	);

	QsysTD_HEX3_HEX0 hex3_hex0 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_hex3_hex0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex3_hex0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex3_hex0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex3_hex0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex3_hex0_s1_readdata),   //                    .readdata
		.out_port   (hex1_export)                                // external_connection.export
	);

	QsysTD_HEX3_HEX0 hex5_hex4 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_hex5_hex4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex5_hex4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex5_hex4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex5_hex4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex5_hex4_s1_readdata),   //                    .readdata
		.out_port   (hex2_export)                                // external_connection.export
	);

	QsysTD_INTERRUPTEURS interrupteurs (
		.clk      (clk_clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address  (mm_interconnect_0_interrupteurs_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_interrupteurs_s1_readdata), //                    .readdata
		.in_port  (interrupteurs_export)                         // external_connection.export
	);

	QsysTD_LEDR ledr (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledr_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	QsysTD_MEMOIRE_ONCHIP memoire_onchip (
		.clk        (clk_clk),                                        //   clk1.clk
		.address    (mm_interconnect_0_memoire_onchip_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memoire_onchip_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memoire_onchip_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memoire_onchip_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memoire_onchip_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memoire_onchip_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memoire_onchip_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	QsysTD_NiosII_CPU niosii_cpu (
		.clk                                 (clk_clk),                                                  //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (niosii_cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (niosii_cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (niosii_cpu_data_master_read),                              //                          .read
		.d_readdata                          (niosii_cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (niosii_cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (niosii_cpu_data_master_write),                             //                          .write
		.d_writedata                         (niosii_cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (niosii_cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (niosii_cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (niosii_cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (niosii_cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (niosii_cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (niosii_cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (niosii_cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (niosii_cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_niosii_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_niosii_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_niosii_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_niosii_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_niosii_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_niosii_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_niosii_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_niosii_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                          // custom_instruction_master.readra
	);

	QsysTD_PWM_CTRL pwm_ctrl (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_pwm_ctrl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pwm_ctrl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pwm_ctrl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pwm_ctrl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pwm_ctrl_s1_readdata),   //                    .readdata
		.out_port   (pwm_ctrl_export)                           // external_connection.export
	);

	QsysTD_PWM_STATUS pwm_status (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_pwm_status_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pwm_status_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pwm_status_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pwm_status_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pwm_status_s1_readdata),   //                    .readdata
		.in_port    (pwm_status_export),                          // external_connection.export
		.irq        (irq_mapper_receiver5_irq)                    //                 irq.irq
	);

	QsysTD_SYS_CLK_timer sys_clk_timer (
		.clk        (clk_clk),                                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               // reset.reset_n
		.address    (mm_interconnect_0_sys_clk_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_clk_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_clk_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_clk_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_clk_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                       //   irq.irq
	);

	QsysTD_SYS_MEL sys_mel (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_sys_mel_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_mel_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_mel_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_mel_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_mel_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                 //   irq.irq
	);

	QsysTD_SYS_SEC sys_sec (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_sys_sec_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_sec_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_sec_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_sec_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_sec_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                 //   irq.irq
	);

	QsysTD_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	QsysTD_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	QsysTD_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                 (clk_clk),                                                     //                               clk_0_clk.clk
		.jtag_uart_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // jtag_uart_0_reset_reset_bridge_in_reset.reset
		.NiosII_CPU_reset_reset_bridge_in_reset_reset  (rst_controller_001_reset_out_reset),                          //  NiosII_CPU_reset_reset_bridge_in_reset.reset
		.NiosII_CPU_data_master_address                (niosii_cpu_data_master_address),                              //                  NiosII_CPU_data_master.address
		.NiosII_CPU_data_master_waitrequest            (niosii_cpu_data_master_waitrequest),                          //                                        .waitrequest
		.NiosII_CPU_data_master_byteenable             (niosii_cpu_data_master_byteenable),                           //                                        .byteenable
		.NiosII_CPU_data_master_read                   (niosii_cpu_data_master_read),                                 //                                        .read
		.NiosII_CPU_data_master_readdata               (niosii_cpu_data_master_readdata),                             //                                        .readdata
		.NiosII_CPU_data_master_write                  (niosii_cpu_data_master_write),                                //                                        .write
		.NiosII_CPU_data_master_writedata              (niosii_cpu_data_master_writedata),                            //                                        .writedata
		.NiosII_CPU_data_master_debugaccess            (niosii_cpu_data_master_debugaccess),                          //                                        .debugaccess
		.NiosII_CPU_instruction_master_address         (niosii_cpu_instruction_master_address),                       //           NiosII_CPU_instruction_master.address
		.NiosII_CPU_instruction_master_waitrequest     (niosii_cpu_instruction_master_waitrequest),                   //                                        .waitrequest
		.NiosII_CPU_instruction_master_read            (niosii_cpu_instruction_master_read),                          //                                        .read
		.NiosII_CPU_instruction_master_readdata        (niosii_cpu_instruction_master_readdata),                      //                                        .readdata
		.NiosII_CPU_instruction_master_readdatavalid   (niosii_cpu_instruction_master_readdatavalid),                 //                                        .readdatavalid
		.BOUTONS_POUSSOIRS_s1_address                  (mm_interconnect_0_boutons_poussoirs_s1_address),              //                    BOUTONS_POUSSOIRS_s1.address
		.BOUTONS_POUSSOIRS_s1_write                    (mm_interconnect_0_boutons_poussoirs_s1_write),                //                                        .write
		.BOUTONS_POUSSOIRS_s1_readdata                 (mm_interconnect_0_boutons_poussoirs_s1_readdata),             //                                        .readdata
		.BOUTONS_POUSSOIRS_s1_writedata                (mm_interconnect_0_boutons_poussoirs_s1_writedata),            //                                        .writedata
		.BOUTONS_POUSSOIRS_s1_chipselect               (mm_interconnect_0_boutons_poussoirs_s1_chipselect),           //                                        .chipselect
		.HEX3_HEX0_s1_address                          (mm_interconnect_0_hex3_hex0_s1_address),                      //                            HEX3_HEX0_s1.address
		.HEX3_HEX0_s1_write                            (mm_interconnect_0_hex3_hex0_s1_write),                        //                                        .write
		.HEX3_HEX0_s1_readdata                         (mm_interconnect_0_hex3_hex0_s1_readdata),                     //                                        .readdata
		.HEX3_HEX0_s1_writedata                        (mm_interconnect_0_hex3_hex0_s1_writedata),                    //                                        .writedata
		.HEX3_HEX0_s1_chipselect                       (mm_interconnect_0_hex3_hex0_s1_chipselect),                   //                                        .chipselect
		.HEX5_HEX4_s1_address                          (mm_interconnect_0_hex5_hex4_s1_address),                      //                            HEX5_HEX4_s1.address
		.HEX5_HEX4_s1_write                            (mm_interconnect_0_hex5_hex4_s1_write),                        //                                        .write
		.HEX5_HEX4_s1_readdata                         (mm_interconnect_0_hex5_hex4_s1_readdata),                     //                                        .readdata
		.HEX5_HEX4_s1_writedata                        (mm_interconnect_0_hex5_hex4_s1_writedata),                    //                                        .writedata
		.HEX5_HEX4_s1_chipselect                       (mm_interconnect_0_hex5_hex4_s1_chipselect),                   //                                        .chipselect
		.INTERRUPTEURS_s1_address                      (mm_interconnect_0_interrupteurs_s1_address),                  //                        INTERRUPTEURS_s1.address
		.INTERRUPTEURS_s1_readdata                     (mm_interconnect_0_interrupteurs_s1_readdata),                 //                                        .readdata
		.jtag_uart_0_avalon_jtag_slave_address         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //           jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                        .write
		.jtag_uart_0_avalon_jtag_slave_read            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                        .read
		.jtag_uart_0_avalon_jtag_slave_readdata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                        .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                        .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                        .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                        .chipselect
		.LEDR_s1_address                               (mm_interconnect_0_ledr_s1_address),                           //                                 LEDR_s1.address
		.LEDR_s1_write                                 (mm_interconnect_0_ledr_s1_write),                             //                                        .write
		.LEDR_s1_readdata                              (mm_interconnect_0_ledr_s1_readdata),                          //                                        .readdata
		.LEDR_s1_writedata                             (mm_interconnect_0_ledr_s1_writedata),                         //                                        .writedata
		.LEDR_s1_chipselect                            (mm_interconnect_0_ledr_s1_chipselect),                        //                                        .chipselect
		.MEMOIRE_ONCHIP_s1_address                     (mm_interconnect_0_memoire_onchip_s1_address),                 //                       MEMOIRE_ONCHIP_s1.address
		.MEMOIRE_ONCHIP_s1_write                       (mm_interconnect_0_memoire_onchip_s1_write),                   //                                        .write
		.MEMOIRE_ONCHIP_s1_readdata                    (mm_interconnect_0_memoire_onchip_s1_readdata),                //                                        .readdata
		.MEMOIRE_ONCHIP_s1_writedata                   (mm_interconnect_0_memoire_onchip_s1_writedata),               //                                        .writedata
		.MEMOIRE_ONCHIP_s1_byteenable                  (mm_interconnect_0_memoire_onchip_s1_byteenable),              //                                        .byteenable
		.MEMOIRE_ONCHIP_s1_chipselect                  (mm_interconnect_0_memoire_onchip_s1_chipselect),              //                                        .chipselect
		.MEMOIRE_ONCHIP_s1_clken                       (mm_interconnect_0_memoire_onchip_s1_clken),                   //                                        .clken
		.NiosII_CPU_debug_mem_slave_address            (mm_interconnect_0_niosii_cpu_debug_mem_slave_address),        //              NiosII_CPU_debug_mem_slave.address
		.NiosII_CPU_debug_mem_slave_write              (mm_interconnect_0_niosii_cpu_debug_mem_slave_write),          //                                        .write
		.NiosII_CPU_debug_mem_slave_read               (mm_interconnect_0_niosii_cpu_debug_mem_slave_read),           //                                        .read
		.NiosII_CPU_debug_mem_slave_readdata           (mm_interconnect_0_niosii_cpu_debug_mem_slave_readdata),       //                                        .readdata
		.NiosII_CPU_debug_mem_slave_writedata          (mm_interconnect_0_niosii_cpu_debug_mem_slave_writedata),      //                                        .writedata
		.NiosII_CPU_debug_mem_slave_byteenable         (mm_interconnect_0_niosii_cpu_debug_mem_slave_byteenable),     //                                        .byteenable
		.NiosII_CPU_debug_mem_slave_waitrequest        (mm_interconnect_0_niosii_cpu_debug_mem_slave_waitrequest),    //                                        .waitrequest
		.NiosII_CPU_debug_mem_slave_debugaccess        (mm_interconnect_0_niosii_cpu_debug_mem_slave_debugaccess),    //                                        .debugaccess
		.PWM_CTRL_s1_address                           (mm_interconnect_0_pwm_ctrl_s1_address),                       //                             PWM_CTRL_s1.address
		.PWM_CTRL_s1_write                             (mm_interconnect_0_pwm_ctrl_s1_write),                         //                                        .write
		.PWM_CTRL_s1_readdata                          (mm_interconnect_0_pwm_ctrl_s1_readdata),                      //                                        .readdata
		.PWM_CTRL_s1_writedata                         (mm_interconnect_0_pwm_ctrl_s1_writedata),                     //                                        .writedata
		.PWM_CTRL_s1_chipselect                        (mm_interconnect_0_pwm_ctrl_s1_chipselect),                    //                                        .chipselect
		.PWM_STATUS_s1_address                         (mm_interconnect_0_pwm_status_s1_address),                     //                           PWM_STATUS_s1.address
		.PWM_STATUS_s1_write                           (mm_interconnect_0_pwm_status_s1_write),                       //                                        .write
		.PWM_STATUS_s1_readdata                        (mm_interconnect_0_pwm_status_s1_readdata),                    //                                        .readdata
		.PWM_STATUS_s1_writedata                       (mm_interconnect_0_pwm_status_s1_writedata),                   //                                        .writedata
		.PWM_STATUS_s1_chipselect                      (mm_interconnect_0_pwm_status_s1_chipselect),                  //                                        .chipselect
		.SYS_CLK_timer_s1_address                      (mm_interconnect_0_sys_clk_timer_s1_address),                  //                        SYS_CLK_timer_s1.address
		.SYS_CLK_timer_s1_write                        (mm_interconnect_0_sys_clk_timer_s1_write),                    //                                        .write
		.SYS_CLK_timer_s1_readdata                     (mm_interconnect_0_sys_clk_timer_s1_readdata),                 //                                        .readdata
		.SYS_CLK_timer_s1_writedata                    (mm_interconnect_0_sys_clk_timer_s1_writedata),                //                                        .writedata
		.SYS_CLK_timer_s1_chipselect                   (mm_interconnect_0_sys_clk_timer_s1_chipselect),               //                                        .chipselect
		.SYS_MEL_s1_address                            (mm_interconnect_0_sys_mel_s1_address),                        //                              SYS_MEL_s1.address
		.SYS_MEL_s1_write                              (mm_interconnect_0_sys_mel_s1_write),                          //                                        .write
		.SYS_MEL_s1_readdata                           (mm_interconnect_0_sys_mel_s1_readdata),                       //                                        .readdata
		.SYS_MEL_s1_writedata                          (mm_interconnect_0_sys_mel_s1_writedata),                      //                                        .writedata
		.SYS_MEL_s1_chipselect                         (mm_interconnect_0_sys_mel_s1_chipselect),                     //                                        .chipselect
		.SYS_SEC_s1_address                            (mm_interconnect_0_sys_sec_s1_address),                        //                              SYS_SEC_s1.address
		.SYS_SEC_s1_write                              (mm_interconnect_0_sys_sec_s1_write),                          //                                        .write
		.SYS_SEC_s1_readdata                           (mm_interconnect_0_sys_sec_s1_readdata),                       //                                        .readdata
		.SYS_SEC_s1_writedata                          (mm_interconnect_0_sys_sec_s1_writedata),                      //                                        .writedata
		.SYS_SEC_s1_chipselect                         (mm_interconnect_0_sys_sec_s1_chipselect),                     //                                        .chipselect
		.sysid_qsys_0_control_slave_address            (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //              sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata           (mm_interconnect_0_sysid_qsys_0_control_slave_readdata)        //                                        .readdata
	);

	QsysTD_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.sender_irq    (niosii_cpu_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (niosii_cpu_debug_reset_request_reset),   // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
